// -------------------------------------------------------------------------
// Portland State University
// Course: ECE585
// 
// Project: L2 Cache Controller
// 
// Filename: L2BUSOP.sv
// 
// Description: Collection of the Bus Operation functions
// -------------------------------------------------------------------------

