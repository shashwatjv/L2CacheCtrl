// -------------------------------------------------------------------------
// Portland State University
// Course: ECE585
// 
// Project: L2 Cache Controller
// 
// Filename: L2CacheCtrl_CfgDefines.svh
// 
// Description: Configuration Defines set to pass parameterized values
// -------------------------------------------------------------------------

`define NUM_PROCESSOR 4
`define PA_BITS 40

`define L1_ASSOC 4
`define L1_LINE_SIZE 32

`define L2_SIZE_KB 16384
`define L2_ASSOC 8
`define L2_LINE_SIZE 64

